module top_module(a,b,c,w,x,y,z);
	input a,b,c;
	output w,x,y,z;
	assign w=a,x=b,y=b,z=c;
endmodule