module top_module(in,out);
	input in;
	output out;
	assign out = in;
endmodule