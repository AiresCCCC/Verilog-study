library verilog;
use verilog.vl_types.all;
entity four_mux_one_tb is
end four_mux_one_tb;
